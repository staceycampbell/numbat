`define RANDOM_CONSTANT 'h54741351
