`define RANDOM_CONSTANT 'h20112C8B
