`define RANDOM_CONSTANT 'h1BD2896C
