`define RANDOM_CONSTANT 1
