module vchess
  (
   input reset,
   input clk
   );

endmodule

