`define RANDOM_CONSTANT 'h38DF46EA
