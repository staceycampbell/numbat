`define WHITE_PAWN 1
`define WHITE_ROOK 2
`define WHITE_KNIT 3
`define WHITE_BISH 4
`define WHITE_KING 5
`define WHITE_QUEN 6

`define BLACK_PAWN 8
`define BLACK_ROOK 9
`define BLACK_KNIT 10
`define BLACK_BISH 11
`define BLACK_KING 12
`define BLACK_QUEN 13

`define PIECE_BITS 4

