`include "vchess.vh"

module vchess_top;

   localparam PIECE_WIDTH = `PIECE_BITS;
   localparam SIDE_WIDTH = PIECE_WIDTH * 8;
   localparam BOARD_WIDTH = PIECE_WIDTH * 8 * 8;
   localparam EVAL_WIDTH = 22;
   localparam MAX_POSITIONS_LOG2 = $clog2(`MAX_POSITIONS);

   integer i;

   reg [BOARD_WIDTH - 1:0] board;
   reg                     board_valid = 0;

   // should be empty
   /*AUTOREGINPUT*/

   /*AUTOWIRE*/
   
   wire                          clk = clk200;

   initial
     begin
        for (i = 0; i < 64; i = i + 1)
          board[i * PIECE_WIDTH+:PIECE_WIDTH] = `EMPTY_POSN;
        board[0 * SIDE_WIDTH + 0 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_ROOK;
        board[0 * SIDE_WIDTH + 1 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_KNIT;
        board[0 * SIDE_WIDTH + 2 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_BISH;
        board[0 * SIDE_WIDTH + 3 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_QUEN;
        board[0 * SIDE_WIDTH + 4 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_KING;
        board[0 * SIDE_WIDTH + 5 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_BISH;
        board[0 * SIDE_WIDTH + 6 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_KNIT;
        board[0 * SIDE_WIDTH + 7 * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_ROOK;
        for (i = 0; i < 8; i = i + 1)
          board[1 * SIDE_WIDTH + i * PIECE_WIDTH+:PIECE_WIDTH] = `WHITE_PAWN;

        board[7 * SIDE_WIDTH + 0 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_ROOK;
        board[7 * SIDE_WIDTH + 1 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_KNIT;
        board[7 * SIDE_WIDTH + 2 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_BISH;
        board[7 * SIDE_WIDTH + 3 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_QUEN;
        board[7 * SIDE_WIDTH + 4 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_KING;
        board[7 * SIDE_WIDTH + 5 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_BISH;
        board[7 * SIDE_WIDTH + 6 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_KNIT;
        board[7 * SIDE_WIDTH + 7 * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_ROOK;
        for (i = 0; i < 8; i = i + 1)
          board[6 * SIDE_WIDTH + i * PIECE_WIDTH+:PIECE_WIDTH] = `BLACK_PAWN;
     end

   always @(posedge clk)
     begin
        board_valid <= 0;
        if (new_board_valid)
          begin
             board <= new_board;
             board_valid <= 1;
          end
     end
   
   /* all_moves AUTO_TEMPLATE (
    .reset (soft_reset),
    .move_count (initial_move_count[]),
    .moves_ready (initial_moves_ready),
    .board_out (initial_board[]),
    .castle_mask_out (initial_castle_mask[]),
    .en_passant_col_out (initial_en_passant_col[]),
    .white_to_move_out (initial_white_to_move),
    .white_in_check_out (initial_white_in_check),
    .black_in_check_out (initial_black_in_check),
    .white_is_attacking_out (initial_white_is_attacking[]),
    .black_is_attacking_out (initial_black_is_attacking[]),
    .capture_out (initial_capture),
    .move_ready (initial_move_ready),
    .\(.*\)_in (\1[]),
    );*/
   all_moves #
     (
      .PIECE_WIDTH (PIECE_WIDTH),
      .SIDE_WIDTH (SIDE_WIDTH),
      .BOARD_WIDTH (BOARD_WIDTH),
      .MAX_POSITIONS_LOG2 (MAX_POSITIONS_LOG2)
      )
   all_moves_initial
     (/*AUTOINST*/
      // Outputs
      .moves_ready                      (initial_moves_ready),   // Templated
      .move_ready                       (initial_move_ready),    // Templated
      .move_count                       (initial_move_count[MAX_POSITIONS_LOG2-1:0]), // Templated
      .board_out                        (initial_board[BOARD_WIDTH-1:0]), // Templated
      .white_to_move_out                (initial_white_to_move), // Templated
      .castle_mask_out                  (initial_castle_mask[3:0]), // Templated
      .en_passant_col_out               (initial_en_passant_col[3:0]), // Templated
      .capture_out                      (initial_capture),       // Templated
      .white_in_check_out               (initial_white_in_check), // Templated
      .black_in_check_out               (initial_black_in_check), // Templated
      .white_is_attacking_out           (initial_white_is_attacking[63:0]), // Templated
      .black_is_attacking_out           (initial_black_is_attacking[63:0]), // Templated
      // Inputs
      .clk                              (clk),
      .reset                            (soft_reset),            // Templated
      .board_valid                      (board_valid),
      .board_in                         (board[BOARD_WIDTH-1:0]), // Templated
      .white_to_move_in                 (white_to_move),         // Templated
      .castle_mask_in                   (castle_mask[3:0]),      // Templated
      .en_passant_col_in                (en_passant_col[3:0]),   // Templated
      .move_index                       (move_index[MAX_POSITIONS_LOG2-1:0]),
      .clear_moves                      (clear_moves));

   reg eval_board_valid;
   reg initial_move_ready_r;

   always @(posedge clk)
     begin
        initial_move_ready_r <= initial_move_ready;
        eval_board_valid <= initial_move_ready && ~initial_move_ready_r;
     end

   /* evaluate AUTO_TEMPLATE (
    .reset (soft_reset),
    .board_in (initial_board[]),
    .board_valid (eval_board_valid),
    .\(.*\)_in (\1[]),
    );*/
   evaluate #
     (
      .PIECE_WIDTH (PIECE_WIDTH),
      .SIDE_WIDTH (SIDE_WIDTH),
      .BOARD_WIDTH (BOARD_WIDTH),
      .EVAL_WIDTH (EVAL_WIDTH)
      )
   evaluate
     (/*AUTOINST*/
      // Outputs
      .eval                             (eval[EVAL_WIDTH-1:0]),
      .eval_valid                       (eval_valid),
      // Inputs
      .clk                              (clk),
      .reset                            (soft_reset),            // Templated
      .board_valid                      (eval_board_valid),      // Templated
      .board_in                         (initial_board[BOARD_WIDTH-1:0]), // Templated
      .white_to_move_in                 (white_to_move),         // Templated
      .castle_mask_in                   (castle_mask[3:0]),      // Templated
      .en_passant_col_in                (en_passant_col[3:0]),   // Templated
      .clear_eval                       (clear_eval));

   /* control AUTO_TEMPLATE (
    );*/
   control #
     (
      .PIECE_WIDTH (PIECE_WIDTH),
      .SIDE_WIDTH (SIDE_WIDTH),
      .BOARD_WIDTH (BOARD_WIDTH),
      .EVAL_WIDTH (EVAL_WIDTH),
      .MAX_POSITIONS_LOG2 (MAX_POSITIONS_LOG2)
      )
   control
     (/*AUTOINST*/
      // Outputs
      .soft_reset                       (soft_reset),
      .new_board                        (new_board[BOARD_WIDTH-1:0]),
      .new_board_valid                  (new_board_valid),
      .castle_mask                      (castle_mask[3:0]),
      .clear_moves                      (clear_moves),
      .en_passant_col                   (en_passant_col[3:0]),
      .white_to_move                    (white_to_move),
      .move_index                       (move_index[MAX_POSITIONS_LOG2-1:0]),
      .clear_eval                       (clear_eval),
      .ctrl0_axi_arready                (ctrl0_axi_arready[0:0]),
      .ctrl0_axi_awready                (ctrl0_axi_awready[0:0]),
      .ctrl0_axi_bresp                  (ctrl0_axi_bresp[1:0]),
      .ctrl0_axi_bvalid                 (ctrl0_axi_bvalid[0:0]),
      .ctrl0_axi_rdata                  (ctrl0_axi_rdata[31:0]),
      .ctrl0_axi_rresp                  (ctrl0_axi_rresp[1:0]),
      .ctrl0_axi_rvalid                 (ctrl0_axi_rvalid[0:0]),
      .ctrl0_axi_wready                 (ctrl0_axi_wready[0:0]),
      .ctrl1_axi_arready                (ctrl1_axi_arready[0:0]),
      .ctrl1_axi_awready                (ctrl1_axi_awready[0:0]),
      .ctrl1_axi_bresp                  (ctrl1_axi_bresp[1:0]),
      .ctrl1_axi_bvalid                 (ctrl1_axi_bvalid[0:0]),
      .ctrl1_axi_rdata                  (ctrl1_axi_rdata[31:0]),
      .ctrl1_axi_rresp                  (ctrl1_axi_rresp[1:0]),
      .ctrl1_axi_rvalid                 (ctrl1_axi_rvalid[0:0]),
      .ctrl1_axi_wready                 (ctrl1_axi_wready[0:0]),
      // Inputs
      .reset                            (reset),
      .clk                              (clk),
      .eval_valid                       (eval_valid),
      .eval                             (eval[EVAL_WIDTH-1:0]),
      .initial_moves_ready              (initial_moves_ready),
      .initial_move_count               (initial_move_count[MAX_POSITIONS_LOG2-1:0]),
      .initial_move_ready               (initial_move_ready),
      .initial_board                    (initial_board[BOARD_WIDTH-1:0]),
      .initial_castle_mask              (initial_castle_mask[3:0]),
      .initial_en_passant_col           (initial_en_passant_col[3:0]),
      .initial_white_to_move            (initial_white_to_move),
      .initial_white_in_check           (initial_white_in_check),
      .initial_black_in_check           (initial_black_in_check),
      .initial_white_is_attacking       (initial_white_is_attacking[63:0]),
      .initial_black_is_attacking       (initial_black_is_attacking[63:0]),
      .initial_capture                  (initial_capture),
      .ctrl0_axi_araddr                 (ctrl0_axi_araddr[39:0]),
      .ctrl0_axi_arprot                 (ctrl0_axi_arprot[2:0]),
      .ctrl0_axi_arvalid                (ctrl0_axi_arvalid),
      .ctrl0_axi_awaddr                 (ctrl0_axi_awaddr[39:0]),
      .ctrl0_axi_awprot                 (ctrl0_axi_awprot[2:0]),
      .ctrl0_axi_awvalid                (ctrl0_axi_awvalid),
      .ctrl0_axi_bready                 (ctrl0_axi_bready),
      .ctrl0_axi_rready                 (ctrl0_axi_rready),
      .ctrl0_axi_wdata                  (ctrl0_axi_wdata[31:0]),
      .ctrl0_axi_wstrb                  (ctrl0_axi_wstrb[3:0]),
      .ctrl0_axi_wvalid                 (ctrl0_axi_wvalid),
      .ctrl1_axi_araddr                 (ctrl1_axi_araddr[39:0]),
      .ctrl1_axi_arprot                 (ctrl1_axi_arprot[2:0]),
      .ctrl1_axi_arvalid                (ctrl1_axi_arvalid),
      .ctrl1_axi_awaddr                 (ctrl1_axi_awaddr[39:0]),
      .ctrl1_axi_awprot                 (ctrl1_axi_awprot[2:0]),
      .ctrl1_axi_awvalid                (ctrl1_axi_awvalid),
      .ctrl1_axi_bready                 (ctrl1_axi_bready),
      .ctrl1_axi_rready                 (ctrl1_axi_rready),
      .ctrl1_axi_wdata                  (ctrl1_axi_wdata[31:0]),
      .ctrl1_axi_wstrb                  (ctrl1_axi_wstrb[3:0]),
      .ctrl1_axi_wvalid                 (ctrl1_axi_wvalid));

   /* mpsoc_preset_wrapper AUTO_TEMPLATE (
    );*/
   mpsoc_preset_wrapper mpsoc_preset_wrapper
     (/*AUTOINST*/);

endmodule

// Local Variables:
// verilog-auto-inst-param-value:t
// verilog-library-directories:(
//     "."
//     "/usr/local/Xilinx/Vivado/2022.1/data/verilog/src/unisims"
//     "vivado/./vchess/vchess_1.gen/sources_1/bd/mpsoc_preset/hdl"
//     )
// End:

