`define EMPTY_POSN (1 << 0)

`define WHITE_PAWN (1 << 1)
`define WHITE_ROOK (1 << 2)
`define WHITE_KNIT (1 << 3)
`define WHITE_BISH (1 << 4)
`define WHITE_KING (1 << 5)
`define WHITE_QUEN (1 << 6)

`define BLACK_PAWN (1 << 8)
`define BLACK_ROOK (1 << 9)
`define BLACK_KNIT (1 << 10)
`define BLACK_BISH (1 << 11)
`define BLACK_KING (1 << 12)
`define BLACK_QUEN (1 << 13)

`define PIECE_BITS 14

`define WHITE_ATTACK 0
`define BLACK_ATTACK 1
